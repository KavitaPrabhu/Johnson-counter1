`timescale 1ns/1ns

// Timing simulation test fixture for jc2_top Verilog design.

module testbench;
   
reg clk;
reg stop;
reg left;
reg right;
wire [3:0] q;
reg PRLD;

jc2_top UUT (
		.left(left),
		.right(right),
		.stop(stop),
		.clk(clk),
		.q(q)
	);

assign glbl.PRLD = PRLD;

initial
begin
	// --------------------
		PRLD = 1;
		clk = 0;
		left = 1;
		right = 1;
		stop = 1;
		// --------------------
		#100
		PRLD = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		left = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		left = 1;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		stop = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		stop = 1;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		right = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		right = 1;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		left = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		left = 1;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;
		// --------------------
		#10
		clk = 1;
		// --------------------
		#10
		clk = 0;

end
endmodule
